// Actuator control electronics
// =============================================================================
// Описание:
// Модуль определитель состояния такотового сигнала.
// =============================================================================

`timescale 1ps / 1ps


/******************************************************************************/
/*-------------------------------- Inclusions --------------------------------*/
/******************************************************************************/
    `include "signals.vh"


/******************************************************************************/
/*---------------------------- Module Description ----------------------------*/
/******************************************************************************/
module CLK_State_Detector_TB
    #(
        parameter TIME_UPDATE_PERIOD_ps = 1000
    )
    (
        input           clk_i,

        output reg[2:0] clk_state_o
    );


/*--------------------------------------------------------------------------*/
/*---------------------------- Local Parameters ----------------------------*/
/*--------------------------------------------------------------------------*/


/******************************************************************************/
/*-------------------------- Signals and  Variables --------------------------*/
/******************************************************************************/
    reg         clk_reg       = 0;
    reg         clk_prev_reg  = 0;


/******************************************************************************/
/*--------------------------------- Behavior ---------------------------------*/
/******************************************************************************/
    /*==================== Main ====================*/
        always #TIME_UPDATE_PERIOD_ps begin
            if (clk_i == clk_prev_reg)
                if (clk_i == 0)
                    clk_state_o = `CLK_STATE_LOW;
                else if (clk_i == 1)
                    clk_state_o = `CLK_STATE_HIGH;
                else
                    clk_state_o = `CLK_STATE_UNDIFINED;
            else if (clk_i != clk_prev_reg)
                if (clk_i == 0)
                    clk_state_o = `CLK_STATE_FALL;
                else if (clk_i == 1)
                    clk_state_o <= `CLK_STATE_RISE;
                else
                    clk_state_o = `CLK_STATE_UNDIFINED;
            else
                clk_state_o = `CLK_STATE_UNDIFINED;
            
            clk_prev_reg = clk_i;
        end
endmodule
