// ////////////////////////////////////////////////////////////////////////////////
// // -*- coding: utf-8; -*-
// // -----------------------------------------------------------------------------
// // [PURPOSE]:   Файл с данными и макросами для работы с числами и математикой.
// //            
// // [FUNCTIONS]: 
// //
// ////////////////////////////////////////////////////////////////////////////////


// `ifndef _math_vh_
//     `define _math_vh_

// /*******************************************************************************/
// /*--------------------------------- Constants ---------------------------------*/
// /*******************************************************************************/
//     /*==================== Math =====================*/
//         `define PI                      3.14159265
//         `define _2PI                    6.283185307


// /*******************************************************************************/
// /*---------------------------- Convertion Factors  ----------------------------*/
// /*******************************************************************************/
//         `define RATIO_DEG_TO_RAD        (2 * `PI / 360)


// `endif