// Actuator control electronics
// ==============================================================================
// Описание:
// Заголовочный файл для работы с модулем SPI.
// ==============================================================================

`ifndef _spi_vh_
    `define _spi_vh_

/*******************************************************************************/
/*-------------------------------- Definitions --------------------------------*/
/*******************************************************************************/
    `define SPI_UPDATE_PERIOD_ps        1000

    `define SPI_ADC_DATA_LEN            12

    /*================= SPI State =================*/
        `define SPI_STATE_IDLE          0
        `define SPI_STATE_TRANSMIT      1
        `define SPI_STATE_SET_RESULT    2
        `define SPI_STATE_FINISH        3
        `define SPI_STATE_ABORT         4


`endif